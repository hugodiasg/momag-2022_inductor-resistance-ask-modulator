** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M_tb-tran.sch
**.subckt ask-915M_tb-tran
Vdd vd GND 3.3
Vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 1500ns 3000ns)
x1 vd out0 in GND ask-915M-0
x2 vd out1 in GND ask-915M-1
x3 vd out2 in GND ask-915M-2
x4 vd out3 in GND ask-915M-3
**** begin user architecture code


*.tran 0.2n 30n
.tran 0.01n 3000n
*.tran 0.3n 400n
*.tran 0.05n 1.3n

.control
destroy all
run

set color0=white
set color1=black
** set hardcopy format
set hcopydevtype=postscript
set hcopypscolor=1

let tol0=maximum(out0)*0.02+0.98*3.3
let tol1=maximum(out1)*0.02+0.98*3.29965
let tol2=maximum(out2)*0.02+0.98*3.29655



plot out0 title 'Out0 - Ideal Inductor'
plot out1 title 'Out1 - R=0.3431 ohms'
plot out2 title 'Out2 - R=3.431 ohms'
plot out3 title 'Out3 - R=34.31 ohms'
plot out0 out1 out2 out3 xlimit 0 10n title 'Out0, Out1, Out2 and Out3'

hardcopy In-915MHz.ps in title 'in - 10MHz'
hardcopy Ideal-915MHz.ps out0 title 'Out0 - Ideal Inductor'
hardcopy Rdiv10-915MHz.ps out1 title 'Out1 - R=0.3431 ohms'
hardcopy R-915MHz.ps out2 title 'Out2 - R=3.431 ohms'
hardcopy Rx10-915MHz.ps out3 title 'Out3 - R=34.31 ohms'
hardcopy Zoom-915MHz.ps out0 out1 out2 out3 xlimit 0 5n title 'Out0, Out1, Out2 and Out3'

*fft out0 out1 out2 out3
*plot mag(out0) mag(out1) mag(out2) mag(out3) xlimit 0.6G 1.6G ylimit 0 7m

*hardcopy fft-915MHz.ps mag(out0) mag(out1) mag(out2) mag(out3) xlimit 0.6G 1.6G ylimit 0 7m

.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-0.sym # of pins=4
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-0.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-0.sch
.subckt ask-915M-0  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=27 L=27 VM=9 m=9
XM1 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
L1 vd out 1.996n m=1
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-1.sym # of pins=4
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-1.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-1.sch
.subckt ask-915M-1  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=27 L=27 VM=9 m=9
XM1 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
x1 vd out l1-915M
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-2.sym # of pins=4
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-2.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-2.sch
.subckt ask-915M-2  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=27 L=27 VM=9 m=9
XM1 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
x1 vd out l2-915M
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-3.sym # of pins=4
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-3.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/ask-915M-3.sch
.subckt ask-915M-3  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=27 L=27 VM=9 m=9
XM1 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
x1 vd out l3-915M
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l1-915M.sym # of pins=2
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l1-915M.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l1-915M.sch
.subckt l1-915M  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.993n m=1
Cs1 p1 net1 147.3f m=1
Cs2 p2 net2 131.8f m=1
Rs1 net1 GND 15.51 m=1
Rs2 net2 GND 8.408 m=1
R1 p2 net3 0.3431 m=1
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l2-915M.sym # of pins=2
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l2-915M.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l2-915M.sch
.subckt l2-915M  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.996n m=1
Cs1 p1 net1 147.3f m=1
Cs2 p2 net2 131.8f m=1
Rs1 net1 GND 15.51 m=1
Rs2 net2 GND 8.408 m=1
R1 p2 net3 3.431 m=1
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l3-915M.sym # of pins=2
** sym_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l3-915M.sym
** sch_path:
*+ /home/hugodg/projects-sky130/sbmo-2022_inductor-resistance-ask-modulator/xschem-915MHz/l3-915M.sch
.subckt l3-915M  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.996n m=1
Cs1 p1 net1 147.3f m=1
Cs2 p2 net2 131.8f m=1
Rs1 net1 GND 15.51 m=1
Rs2 net2 GND 8.408 m=1
R1 p2 net3 34.31 m=1
.ends

.GLOBAL GND
.end
